-- Copyright (C) 2022  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 21.1.1 Build 850 06/23/2022 SJ Lite Edition"
-- CREATED		"Sun Nov 13 23:02:46 2022"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY f4b IS 
	PORT
	(
		clk :  IN  STD_LOGIC;
		reset :  IN  STD_LOGIC;
		clkMBR :  IN  STD_LOGIC;
		ACC :  OUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		BR_OUT :  OUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		BRIN :  OUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		CAROUT :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0);
		CONTROL :  OUT  STD_LOGIC_VECTOR(31 DOWNTO 0);
		IROUT :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0);
		MAROUT :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0);
		PC :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0);
		RAM_OUT :  OUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		RAMIN :  OUT  STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END f4b;

ARCHITECTURE bdf_type OF f4b IS 

ATTRIBUTE black_box : BOOLEAN;
ATTRIBUTE noopt : BOOLEAN;

COMPONENT lpm_ram_dq_1
	PORT(inclock : IN STD_LOGIC;
		 we : IN STD_LOGIC;
		 address : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 data : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_ram_dq_1: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_ram_dq_1: COMPONENT IS true;

COMPONENT lpm_rom_0
	PORT(inclock : IN STD_LOGIC;
		 address : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(31 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF lpm_rom_0: COMPONENT IS true;
ATTRIBUTE noopt OF lpm_rom_0: COMPONENT IS true;

COMPONENT alu
	PORT(clk : IN STD_LOGIC;
		 reset : IN STD_LOGIC;
		 ACCclear : IN STD_LOGIC;
		 aluCONTR : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 BR : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 PCjmp : OUT STD_LOGIC;
		 ACC : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT br
	PORT(MBR_BRc : IN STD_LOGIC;
		 MBR_BR : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 BRout : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT car
	PORT(clk : IN STD_LOGIC;
		 reset : IN STD_LOGIC;
		 CAR : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 CARc : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 OP : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 CARout : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT controlr
	PORT(control : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 R : OUT STD_LOGIC;
		 W : OUT STD_LOGIC;
		 RW : OUT STD_LOGIC;
		 PCc1 : OUT STD_LOGIC;
		 PCinc : OUT STD_LOGIC;
		 PCc3 : OUT STD_LOGIC;
		 ACCclear : OUT STD_LOGIC;
		 MBR_MARc : OUT STD_LOGIC;
		 PC_MARc : OUT STD_LOGIC;
		 ACC_MBRc : OUT STD_LOGIC;
		 MBR_OPc : OUT STD_LOGIC;
		 MBR_BRc : OUT STD_LOGIC;
		 CAR : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 CARc : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 CONTRout : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

COMPONENT ir
	PORT(opcode : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 IRout : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT mar
	PORT(clk : IN STD_LOGIC;
		 PC_MARc : IN STD_LOGIC;
		 MBR_MARc : IN STD_LOGIC;
		 MBR_MAR : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 PC : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 MARout : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT mbr
	PORT(clk : IN STD_LOGIC;
		 reset : IN STD_LOGIC;
		 MBR_OPc : IN STD_LOGIC;
		 ACC_MBRc : IN STD_LOGIC;
		 R : IN STD_LOGIC;
		 W : IN STD_LOGIC;
		 ACC_MBR : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 RAM_MBR : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 MBR_BR : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 MBR_MAR : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 MBR_OP : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 MBR_PC : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 MBR_RAM : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT pc
	PORT(clk : IN STD_LOGIC;
		 PCjmp : IN STD_LOGIC;
		 PCc1 : IN STD_LOGIC;
		 PCinc : IN STD_LOGIC;
		 PCc3 : IN STD_LOGIC;
		 reset : IN STD_LOGIC;
		 CONTRalu : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 MBR_PC : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 PCout : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC_VECTOR(7 DOWNTO 0);


BEGIN 
ACC <= SYNTHESIZED_WIRE_22;
BR_OUT <= SYNTHESIZED_WIRE_2;
BRIN <= SYNTHESIZED_WIRE_8;
CAROUT <= SYNTHESIZED_WIRE_3;
CONTROL <= SYNTHESIZED_WIRE_12;
IROUT <= SYNTHESIZED_WIRE_11;
MAROUT <= SYNTHESIZED_WIRE_5;
PC <= SYNTHESIZED_WIRE_17;
RAM_OUT <= SYNTHESIZED_WIRE_23;
RAMIN <= SYNTHESIZED_WIRE_6;



b2v_inst : alu
PORT MAP(clk => clk,
		 reset => reset,
		 ACCclear => SYNTHESIZED_WIRE_0,
		 aluCONTR => SYNTHESIZED_WIRE_30,
		 BR => SYNTHESIZED_WIRE_2,
		 PCjmp => SYNTHESIZED_WIRE_24,
		 ACC => SYNTHESIZED_WIRE_22);


b2v_inst13 : lpm_rom_0
PORT MAP(inclock => clk,
		 address => SYNTHESIZED_WIRE_3,
		 q => SYNTHESIZED_WIRE_12);


b2v_inst14 : lpm_ram_dq_1
PORT MAP(inclock => clk,
		 we => SYNTHESIZED_WIRE_4,
		 address => SYNTHESIZED_WIRE_5,
		 data => SYNTHESIZED_WIRE_6,
		 q => SYNTHESIZED_WIRE_23);


b2v_inst2 : br
PORT MAP(MBR_BRc => SYNTHESIZED_WIRE_7,
		 MBR_BR => SYNTHESIZED_WIRE_8,
		 BRout => SYNTHESIZED_WIRE_2);


b2v_inst3 : car
PORT MAP(clk => clk,
		 reset => reset,
		 CAR => SYNTHESIZED_WIRE_9,
		 CARc => SYNTHESIZED_WIRE_10,
		 OP => SYNTHESIZED_WIRE_11,
		 CARout => SYNTHESIZED_WIRE_3);


b2v_inst4 : controlr
PORT MAP(control => SYNTHESIZED_WIRE_12,
		 R => SYNTHESIZED_WIRE_20,
		 W => SYNTHESIZED_WIRE_21,
		 RW => SYNTHESIZED_WIRE_4,
		 PCc1 => SYNTHESIZED_WIRE_25,
		 PCinc => SYNTHESIZED_WIRE_26,
		 PCc3 => SYNTHESIZED_WIRE_27,
		 ACCclear => SYNTHESIZED_WIRE_0,
		 MBR_MARc => SYNTHESIZED_WIRE_15,
		 PC_MARc => SYNTHESIZED_WIRE_14,
		 ACC_MBRc => SYNTHESIZED_WIRE_19,
		 MBR_OPc => SYNTHESIZED_WIRE_18,
		 MBR_BRc => SYNTHESIZED_WIRE_7,
		 CAR => SYNTHESIZED_WIRE_9,
		 CARc => SYNTHESIZED_WIRE_10,
		 CONTRout => SYNTHESIZED_WIRE_30);


b2v_inst5 : ir
PORT MAP(opcode => SYNTHESIZED_WIRE_13,
		 IRout => SYNTHESIZED_WIRE_11);


b2v_inst6 : mar
PORT MAP(clk => clk,
		 PC_MARc => SYNTHESIZED_WIRE_14,
		 MBR_MARc => SYNTHESIZED_WIRE_15,
		 MBR_MAR => SYNTHESIZED_WIRE_16,
		 PC => SYNTHESIZED_WIRE_17,
		 MARout => SYNTHESIZED_WIRE_5);


b2v_inst7 : mbr
PORT MAP(clk => clkMBR,
		 reset => reset,
		 MBR_OPc => SYNTHESIZED_WIRE_18,
		 ACC_MBRc => SYNTHESIZED_WIRE_19,
		 R => SYNTHESIZED_WIRE_20,
		 W => SYNTHESIZED_WIRE_21,
		 ACC_MBR => SYNTHESIZED_WIRE_22,
		 RAM_MBR => SYNTHESIZED_WIRE_23,
		 MBR_BR => SYNTHESIZED_WIRE_8,
		 MBR_MAR => SYNTHESIZED_WIRE_16,
		 MBR_OP => SYNTHESIZED_WIRE_13,
		 MBR_PC => SYNTHESIZED_WIRE_29,
		 MBR_RAM => SYNTHESIZED_WIRE_6);


b2v_inst8 : pc
PORT MAP(clk => clk,
		 PCjmp => SYNTHESIZED_WIRE_24,
		 PCc1 => SYNTHESIZED_WIRE_25,
		 PCinc => SYNTHESIZED_WIRE_26,
		 PCc3 => SYNTHESIZED_WIRE_27,
		 reset => reset,
		 CONTRalu => SYNTHESIZED_WIRE_30,
		 MBR_PC => SYNTHESIZED_WIRE_29,
		 PCout => SYNTHESIZED_WIRE_17);


END bdf_type;